* NGSPICE file created from CLS.ext - technology: sky130A

.subckt CLS VIN VDDH VOUT GND VDDL
X0 A VIN GND GND sky130_fd_pr__nfet_01v8 ad=0.246 pd=2.02 as=0.234 ps=1.98 w=0.6 l=0.2
X1 A VIN VDDL VDDL sky130_fd_pr__pfet_01v8 ad=0.246 pd=2.02 as=0.234 ps=1.98 w=0.6 l=0.2
X2 a_250_n620# E VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=2 pd=9 as=1.6 ps=4.8 w=4 l=0.8
X3 VOUT E VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=3 pd=11.2 as=3 ps=11.2 w=5 l=0.5
X4 a_180_n1399# A GND GND sky130_fd_pr__nfet_01v8 ad=1.2 pd=8.6 as=1.2 ps=4.6 w=4 l=0.15
X5 VOUT E GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.2 pd=5.2 as=1.2 ps=5.2 w=2 l=0.5
X6 GND VIN a_60_n1399# GND sky130_fd_pr__nfet_01v8 ad=1.2 pd=4.6 as=1.2 ps=8.6 w=4 l=0.15
X7 VDDH G a_n40_n620# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=1.6 pd=4.8 as=2 ps=9 w=4 l=0.8
.ends

