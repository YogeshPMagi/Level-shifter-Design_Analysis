magic
tech sky130A
timestamp 1771746969
<< nwell >>
rect -80 -655 550 -80
rect 306 -754 550 -655
rect -230 -1178 -90 -1020
<< nmos >>
rect -170 -1287 -150 -1227
rect 90 -1399 105 -999
rect 165 -1399 180 -999
<< pmos >>
rect -170 -1160 -150 -1100
<< mvnmos >>
rect 400 -1060 450 -860
<< mvpmos >>
rect 10 -620 90 -220
rect 170 -620 250 -220
rect 400 -720 450 -220
<< ndiff >>
rect 60 -1007 90 -999
rect -209 -1235 -170 -1227
rect -209 -1279 -201 -1235
rect -177 -1279 -170 -1235
rect -209 -1287 -170 -1279
rect -150 -1235 -109 -1227
rect -150 -1279 -141 -1235
rect -117 -1279 -109 -1235
rect -150 -1287 -109 -1279
rect 60 -1391 65 -1007
rect 82 -1391 90 -1007
rect 60 -1399 90 -1391
rect 105 -1007 165 -999
rect 105 -1391 111 -1007
rect 159 -1391 165 -1007
rect 105 -1399 165 -1391
rect 180 -1007 210 -999
rect 180 -1391 188 -1007
rect 205 -1391 210 -1007
rect 180 -1399 210 -1391
<< pdiff >>
rect -209 -1108 -170 -1100
rect -209 -1152 -201 -1108
rect -177 -1152 -170 -1108
rect -209 -1160 -170 -1152
rect -150 -1108 -109 -1100
rect -150 -1152 -141 -1108
rect -117 -1152 -109 -1108
rect -150 -1160 -109 -1152
<< mvndiff >>
rect 340 -870 400 -860
rect 340 -1050 350 -870
rect 390 -1050 400 -870
rect 340 -1060 400 -1050
rect 450 -870 510 -860
rect 450 -1050 460 -870
rect 500 -1050 510 -870
rect 450 -1060 510 -1050
<< mvpdiff >>
rect -40 -230 10 -220
rect -40 -610 -30 -230
rect 0 -610 10 -230
rect -40 -620 10 -610
rect 90 -230 170 -220
rect 90 -610 100 -230
rect 160 -610 170 -230
rect 90 -620 170 -610
rect 250 -230 300 -220
rect 250 -610 259 -230
rect 290 -610 300 -230
rect 250 -620 300 -610
rect 340 -230 400 -220
rect 340 -710 350 -230
rect 390 -710 400 -230
rect 340 -720 400 -710
rect 450 -230 510 -220
rect 450 -710 460 -230
rect 500 -710 510 -230
rect 450 -720 510 -710
<< ndiffc >>
rect -201 -1279 -177 -1235
rect -141 -1279 -117 -1235
rect 65 -1391 82 -1007
rect 111 -1391 159 -1007
rect 188 -1391 205 -1007
<< pdiffc >>
rect -201 -1152 -177 -1108
rect -141 -1152 -117 -1108
<< mvndiffc >>
rect 350 -1050 390 -870
rect 460 -1050 500 -870
<< mvpdiffc >>
rect -30 -610 0 -230
rect 100 -610 160 -230
rect 259 -610 290 -230
rect 350 -710 390 -230
rect 460 -710 500 -230
<< psubdiff >>
rect -210 -1322 -107 -1314
rect -210 -1342 -198 -1322
rect -120 -1342 -107 -1322
rect -210 -1349 -107 -1342
<< nsubdiff >>
rect -211 -1046 -108 -1038
rect -211 -1066 -198 -1046
rect -120 -1066 -108 -1046
rect -211 -1073 -108 -1066
<< mvpsubdiff >>
rect 335 -1143 496 -1132
rect 335 -1160 348 -1143
rect 482 -1160 496 -1143
rect 335 -1168 496 -1160
rect -40 -1455 300 -1446
rect -40 -1478 -27 -1455
rect 287 -1478 300 -1455
rect -40 -1487 300 -1478
<< mvnsubdiff >>
rect -40 -128 510 -121
rect -40 -151 -27 -128
rect 287 -151 340 -128
rect -40 -152 340 -151
rect 485 -152 510 -128
rect -40 -160 510 -152
rect -40 -161 299 -160
<< psubdiffcont >>
rect -198 -1342 -120 -1322
<< nsubdiffcont >>
rect -198 -1066 -120 -1046
<< mvpsubdiffcont >>
rect 348 -1160 482 -1143
rect -27 -1478 287 -1455
<< mvnsubdiffcont >>
rect -27 -151 287 -128
rect 340 -152 485 -128
<< poly >>
rect 10 -220 90 -207
rect 170 -220 250 -207
rect 400 -220 450 -207
rect 10 -667 90 -620
rect 10 -677 108 -667
rect 10 -737 32 -677
rect 98 -737 108 -677
rect 10 -747 108 -737
rect 170 -761 250 -620
rect 151 -771 250 -761
rect 151 -831 161 -771
rect 227 -831 250 -771
rect 151 -841 250 -831
rect 400 -770 450 -720
rect 400 -830 410 -770
rect 440 -830 450 -770
rect 400 -860 450 -830
rect 81 -901 115 -896
rect 81 -921 90 -901
rect 107 -921 115 -901
rect 81 -926 115 -921
rect 90 -999 105 -926
rect 155 -957 189 -952
rect 155 -977 164 -957
rect 181 -977 189 -957
rect 155 -982 189 -977
rect 165 -999 180 -982
rect -170 -1100 -150 -1087
rect -170 -1179 -150 -1160
rect -191 -1185 -150 -1179
rect -191 -1202 -183 -1185
rect -166 -1202 -150 -1185
rect -191 -1210 -150 -1202
rect -170 -1227 -150 -1210
rect -170 -1300 -150 -1287
rect 400 -1073 450 -1060
rect 90 -1412 105 -1399
rect 165 -1412 180 -1399
<< polycont >>
rect 32 -737 98 -677
rect 161 -831 227 -771
rect 410 -830 440 -770
rect 90 -921 107 -901
rect 164 -977 181 -957
rect -183 -1202 -166 -1185
<< locali >>
rect -40 -128 100 -121
rect 160 -128 510 -121
rect -40 -151 -27 -128
rect 287 -151 340 -128
rect -40 -161 100 -151
rect 160 -152 340 -151
rect 485 -152 510 -128
rect 160 -160 510 -152
rect 160 -161 299 -160
rect -40 -230 9 -220
rect -40 -400 -30 -230
rect -40 -430 -32 -400
rect -40 -610 -30 -430
rect 0 -610 9 -230
rect -40 -620 9 -610
rect 90 -230 169 -220
rect 90 -610 100 -230
rect 160 -610 169 -230
rect 90 -620 169 -610
rect 250 -230 300 -220
rect 250 -610 259 -230
rect 290 -400 300 -230
rect 291 -430 300 -400
rect 290 -610 300 -430
rect 250 -620 300 -610
rect 340 -230 400 -220
rect 23 -677 108 -667
rect 23 -737 32 -677
rect 98 -737 108 -677
rect 340 -710 350 -230
rect 390 -710 400 -230
rect 340 -720 400 -710
rect 450 -230 510 -220
rect 450 -710 460 -230
rect 500 -710 510 -230
rect 450 -720 510 -710
rect 23 -747 108 -737
rect 151 -771 236 -761
rect 151 -831 161 -771
rect 227 -831 236 -771
rect 151 -841 236 -831
rect 400 -770 450 -761
rect 400 -830 410 -770
rect 440 -830 450 -770
rect 400 -841 450 -830
rect 340 -870 400 -860
rect 81 -901 115 -896
rect 81 -921 90 -901
rect 107 -921 115 -901
rect 81 -926 115 -921
rect 155 -957 189 -952
rect 155 -977 164 -957
rect 181 -977 189 -957
rect 155 -982 189 -977
rect 60 -1007 90 -999
rect -211 -1046 -108 -1038
rect -211 -1047 -198 -1046
rect -211 -1065 -201 -1047
rect -211 -1066 -198 -1065
rect -120 -1066 -108 -1046
rect -211 -1073 -108 -1066
rect -201 -1100 -177 -1073
rect -209 -1108 -170 -1100
rect -209 -1152 -201 -1108
rect -177 -1152 -170 -1108
rect -209 -1160 -170 -1152
rect -150 -1108 -109 -1100
rect -150 -1152 -141 -1108
rect -117 -1152 -109 -1108
rect -150 -1160 -109 -1152
rect -191 -1185 -158 -1179
rect -191 -1202 -183 -1185
rect -166 -1202 -158 -1185
rect -191 -1210 -158 -1202
rect -141 -1183 -117 -1160
rect -141 -1206 -135 -1183
rect -141 -1227 -117 -1206
rect -209 -1235 -170 -1227
rect -209 -1279 -201 -1235
rect -177 -1279 -170 -1235
rect -209 -1287 -170 -1279
rect -150 -1235 -109 -1227
rect -150 -1279 -141 -1235
rect -117 -1279 -109 -1235
rect -150 -1287 -109 -1279
rect -201 -1314 -177 -1287
rect -210 -1322 -107 -1314
rect -210 -1323 -198 -1322
rect -210 -1341 -200 -1323
rect -210 -1342 -198 -1341
rect -120 -1342 -107 -1322
rect -210 -1349 -107 -1342
rect 60 -1391 65 -1007
rect 82 -1391 90 -1007
rect 60 -1399 90 -1391
rect 107 -1007 163 -999
rect 107 -1391 111 -1007
rect 159 -1391 163 -1007
rect 107 -1399 163 -1391
rect 180 -1007 210 -999
rect 180 -1391 188 -1007
rect 205 -1391 210 -1007
rect 340 -1050 350 -870
rect 390 -1050 400 -870
rect 340 -1060 400 -1050
rect 450 -870 510 -860
rect 450 -1050 460 -870
rect 500 -1050 510 -870
rect 450 -1060 510 -1050
rect 350 -1132 390 -1130
rect 335 -1143 496 -1132
rect 335 -1160 348 -1143
rect 482 -1160 496 -1143
rect 335 -1168 496 -1160
rect 180 -1399 210 -1391
rect 111 -1446 159 -1399
rect -40 -1449 300 -1446
rect -40 -1455 100 -1449
rect 170 -1455 300 -1449
rect -40 -1478 -27 -1455
rect 287 -1478 300 -1455
rect -40 -1483 100 -1478
rect 170 -1483 300 -1478
rect -40 -1487 300 -1483
<< viali >>
rect 100 -128 160 -120
rect 100 -151 160 -128
rect 100 -160 160 -151
rect 350 -152 390 -128
rect -32 -430 -30 -400
rect -30 -430 0 -400
rect 104 -430 156 -400
rect 259 -430 290 -400
rect 290 -430 291 -400
rect 32 -737 98 -677
rect 353 -480 387 -450
rect 463 -480 497 -450
rect 161 -831 227 -771
rect 410 -830 440 -770
rect 90 -921 107 -901
rect 164 -977 181 -957
rect -201 -1065 -198 -1047
rect -198 -1065 -177 -1047
rect -183 -1202 -166 -1185
rect -135 -1206 -114 -1183
rect -200 -1341 -198 -1323
rect -198 -1341 -178 -1323
rect 65 -1210 82 -1180
rect 188 -1210 205 -1180
rect 353 -970 387 -950
rect 463 -970 497 -950
rect 350 -1160 390 -1143
rect 100 -1455 170 -1449
rect 100 -1478 170 -1455
rect 100 -1483 170 -1478
<< metal1 >>
rect -60 -110 533 -109
rect -120 -120 589 -110
rect -120 -160 100 -120
rect 160 -128 589 -120
rect 160 -152 350 -128
rect 390 -152 589 -128
rect 160 -160 589 -152
rect -120 -170 589 -160
rect -40 -400 10 -370
rect -40 -430 -32 -400
rect 0 -430 10 -400
rect -40 -431 10 -430
rect 100 -400 160 -170
rect 100 -430 104 -400
rect 156 -430 160 -400
rect -40 -766 9 -431
rect 100 -460 160 -430
rect 250 -400 300 -370
rect 250 -430 259 -400
rect 291 -430 300 -400
rect 23 -677 109 -667
rect 23 -737 32 -677
rect 99 -737 109 -677
rect 23 -747 109 -737
rect 250 -673 300 -430
rect 350 -450 390 -170
rect 350 -480 353 -450
rect 387 -480 390 -450
rect 350 -510 390 -480
rect 460 -450 500 -430
rect 460 -480 463 -450
rect 497 -480 500 -450
rect 250 -743 255 -673
rect 296 -743 300 -673
rect 250 -748 300 -743
rect -40 -837 -36 -766
rect 6 -837 9 -766
rect -40 -841 9 -837
rect 150 -766 236 -761
rect 150 -836 156 -766
rect 230 -836 236 -766
rect 150 -841 236 -836
rect -40 -1000 -10 -841
rect 81 -898 115 -896
rect 81 -924 84 -898
rect 112 -924 115 -898
rect 81 -926 115 -924
rect 155 -954 189 -952
rect 155 -980 158 -954
rect 186 -980 189 -954
rect 155 -982 189 -980
rect 180 -1000 210 -999
rect 270 -1000 300 -748
rect 404 -770 446 -764
rect 404 -831 410 -770
rect 440 -831 446 -770
rect 404 -837 446 -831
rect 460 -770 500 -480
rect 460 -831 470 -770
rect 497 -831 500 -770
rect -40 -1030 90 -1000
rect -225 -1047 -95 -1038
rect -225 -1065 -201 -1047
rect -177 -1065 -95 -1047
rect -225 -1073 -95 -1065
rect -191 -1181 -158 -1179
rect -191 -1208 -188 -1181
rect -161 -1208 -158 -1181
rect -191 -1210 -158 -1208
rect -141 -1180 -108 -1179
rect -141 -1209 -138 -1180
rect -111 -1209 -108 -1180
rect -141 -1210 -108 -1209
rect 60 -1180 90 -1030
rect 60 -1210 65 -1180
rect 82 -1210 90 -1180
rect 180 -1029 300 -1000
rect 350 -950 390 -860
rect 350 -970 353 -950
rect 387 -970 390 -950
rect 180 -1180 210 -1029
rect 350 -1130 390 -970
rect 460 -950 500 -831
rect 460 -970 463 -950
rect 497 -970 500 -950
rect 460 -1060 500 -970
rect 330 -1143 500 -1130
rect 330 -1160 350 -1143
rect 390 -1160 500 -1143
rect 330 -1170 500 -1160
rect 60 -1260 90 -1210
rect -222 -1323 -92 -1314
rect -222 -1341 -200 -1323
rect -178 -1341 -92 -1323
rect -222 -1349 -92 -1341
rect 111 -1440 159 -1195
rect 180 -1210 188 -1180
rect 205 -1210 210 -1180
rect 180 -1260 210 -1210
rect -50 -1449 310 -1440
rect -50 -1483 100 -1449
rect 170 -1483 310 -1449
rect -50 -1490 310 -1483
<< via1 >>
rect 32 -737 98 -677
rect 98 -737 99 -677
rect 255 -743 296 -673
rect -36 -837 6 -766
rect 156 -771 230 -766
rect 156 -831 161 -771
rect 161 -831 227 -771
rect 227 -831 230 -771
rect 156 -836 230 -831
rect 84 -901 112 -898
rect 84 -921 90 -901
rect 90 -921 107 -901
rect 107 -921 112 -901
rect 84 -924 112 -921
rect 158 -957 186 -954
rect 158 -977 164 -957
rect 164 -977 181 -957
rect 181 -977 186 -957
rect 158 -980 186 -977
rect 410 -830 440 -770
rect 410 -831 440 -830
rect 470 -831 497 -770
rect -188 -1185 -161 -1181
rect -188 -1202 -183 -1185
rect -183 -1202 -166 -1185
rect -166 -1202 -161 -1185
rect -188 -1208 -161 -1202
rect -138 -1183 -111 -1180
rect -138 -1206 -135 -1183
rect -135 -1206 -114 -1183
rect -114 -1206 -111 -1183
rect -138 -1209 -111 -1206
<< metal2 >>
rect 23 -673 300 -667
rect 23 -677 255 -673
rect 23 -737 32 -677
rect 99 -737 255 -677
rect 23 -743 255 -737
rect 296 -743 300 -673
rect 23 -747 300 -743
rect -40 -766 450 -761
rect -40 -837 -36 -766
rect 6 -836 156 -766
rect 230 -770 450 -766
rect 230 -831 410 -770
rect 440 -831 450 -770
rect 230 -836 450 -831
rect 6 -837 450 -836
rect -40 -841 450 -837
rect 467 -770 683 -760
rect 467 -831 470 -770
rect 497 -831 683 -770
rect 467 -840 683 -831
rect -265 -905 -250 -865
rect 81 -898 115 -896
rect 81 -905 84 -898
rect -265 -920 84 -905
rect -265 -1185 -250 -920
rect 81 -924 84 -920
rect 112 -924 115 -898
rect 81 -926 115 -924
rect 155 -954 189 -952
rect 155 -960 158 -954
rect -70 -975 158 -960
rect -191 -1181 -158 -1179
rect -191 -1185 -188 -1181
rect -265 -1200 -188 -1185
rect -191 -1208 -188 -1200
rect -161 -1208 -158 -1181
rect -191 -1210 -158 -1208
rect -141 -1180 -108 -1179
rect -141 -1209 -138 -1180
rect -111 -1185 -108 -1180
rect -70 -1185 -55 -975
rect 155 -980 158 -975
rect 186 -980 189 -954
rect 155 -982 189 -980
rect -111 -1200 -55 -1185
rect -111 -1209 -108 -1200
rect -141 -1210 -108 -1209
<< labels >>
rlabel metal1 537 -140 537 -140 1 VDDH
port 2 n default bidirectional
rlabel metal1 -214 -1344 -214 -1344 1 GND
port 4 n default bidirectional
rlabel metal1 -37 -1468 -37 -1468 1 GND
port 4 n default bidirectional
rlabel metal1 338 -1153 338 -1153 1 GND
port 4 n default bidirectional
rlabel metal2 -111 -1200 -55 -1185 1 A
rlabel metal2 -70 -975 158 -960 1 A
rlabel metal2 -259 -889 -256 -868 1 VIN
port 1 n default input
rlabel metal1 460 -1060 467 -470 1 F
rlabel metal1 245 -1011 245 -1011 1 G
rlabel metal1 6 -1011 6 -1011 1 H
rlabel metal2 141 -702 141 -702 1 I
rlabel space 59 -1399 89 -999 1 N
rlabel nwell -40 -620 10 -220 1 O
rlabel metal2 570 -803 594 -797 1 VOUT
port 3 n default output
rlabel metal2 609 -796 609 -796 1 VOUT
port 3 n default output
rlabel metal1 -205 -1058 -202 -1054 1 VDDL
port 5 n
rlabel metal1 250 -620 300 -370 1 M
rlabel metal1 100 -170 160 -160 1 B
rlabel metal1 350 -230 390 -152 1 C
rlabel metal1 60 -1399 90 -1349 1 K
<< end >>
