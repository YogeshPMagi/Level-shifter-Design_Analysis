** sch_path: /home/yogesh/   DCVSL.sch
**.subckt    DCVSL
XMp3 net1 o VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 L=0.80 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMp4 VOUT o VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 L=0.50 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMN4 VOUT o GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.50 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
VIN VIN GND pulse(0 1.2 1n 0.3n 0.3n 5n 10n)
VSS1 VDDH GND 3.3v
XMN2 o VIN GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
VDD VDDl GND 1.2v
XMN3 net1 i GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMp2 o net1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 L=0.80 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMN1 i VIN GND GND sky130_fd_pr__nfet_01v8 L=0.2 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMP1 i VIN VDDl VDDl sky130_fd_pr__pfet_01v8 L=0.2 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code


.lib /home/yogesh/OpenLane/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
* Perfect Timing Analysis
.tran 0.01n 50n
* Measure 10% to 90% Rise Time (The slope going up)
.meas tran rise_time trig v(vout) val=0.33 rise=1 targ v(vout) val=2.97 rise=1
* Measure 90% to 10% Fall Time (The slope going down)
.meas tran fall_time trig v(vout) val=2.97 fall=1 targ v(vout) val=0.33 fall=1
* 1. Timing Measurements (50% to 50% for Prop Delay)
.meas tran t_plh trig v(vin) val=0.6 rise=1 targ v(vout) val=1.65 rise=1
.meas tran t_phl trig v(vin) val=0.6 fall=1 targ v(vout) val=1.65 fall=1
.meas tran energy_total integ vss1#branch

**** end user architecture code
**.ends
.GLOBAL GND
.end
